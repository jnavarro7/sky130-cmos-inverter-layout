* SPICE3 file created from inverter.ext - technology: sky130A

.option scale=10m

X0 a_15_n15# a_n25_n75# a_n65_n15# w_n90_n40# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0 l=0
X1 a_15_n140# a_n25_n75# a_n50_n140# SUB sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0 l=0
